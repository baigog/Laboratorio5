library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY RS232_FSM IS
	PORT(
	DATA_READY: IN STD_LOGIC;
	SR_DONE:		IN	STD_LOGIC;
	CLK:			IN STD_LOGIC;
	RST:			IN	STD_LOGIC;
	
	BUSY:			OUT	STD_LOGIC;
	SHIFT:		OUT	STD_LOGIC;
	SS:			OUT	STD_LOGIC;
	SEL:			OUT	STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END RS232_FSM;

ARCHITECTURE BEH OF RS232_FSM IS
TYPE STATE IS (INIT,IDLE,START,DATA,PARITY);
SIGNAL CS,NS: STATE;

BEGIN

NEXT_STATE: PROCESS (CS,DATA_READY,SR_DONE)
BEGIN
	CASE CS IS
		WHEN IDLE	=>
			IF	(DATA_READY='1')	THEN
				NS	<=	START;
			ELSE
				NS	<=	IDLE;
			END IF;
		WHEN START	=>
			NS<= DATA;
		WHEN DATA	=>
			IF	(SR_DONE='1')	THEN
				NS	<=	PARITY;
			ELSE
				NS <=	DATA;
			END IF;
		WHEN PARITY	=>
			NS	<=	IDLE;
		WHEN OTHERS	=>
			NS	<=	IDLE;
	END CASE;
END PROCESS;

CURRENT_STATE: PROCESS (CLK, RST)
BEGIN
	IF	(RST='1') THEN
		CS <= IDLE;
	ELSIF	(RISING_EDGE(CLK)) THEN
		CS <= NS;
	END IF;
END PROCESS;

OUTPUTS:	PROCESS (CLK,RST)
BEGIN
	IF	(RST='1') THEN
		SHIFT<='0';
		SS<='1';
		SEL<="00";
		BUSY<='0';
	ELSIF(RISING_EDGE(CLK)) THEN
		BUSY<='1';
		SHIFT<='0';
		SS<='1';
		SEL<="00";
		CASE CS IS
			WHEN IDLE	=> BUSY<='0';
			WHEN START	=>
				SS<='0';
			WHEN DATA	=>
				SEL<="01";
				SHIFT<='1';
			WHEN PARITY	=>
				SEL<="11";
			WHEN OTHERS	=> NULL;
		END CASE;
	END IF;
END PROCESS;
END BEH;
	 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
ENTITY SHIFT_REGISTER IS
PORT(
	CLK:				IN		STD_LOGIC;
	RST:				IN		STD_LOGIC;
	DATAIN:			IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
	SHIFT_LOAD:		IN		STD_LOGIC_VECTOR(1 DOWNTO 0);	--01: SHIFT	1X: LOAD	00: DO NOTHING
	DATAOUT:			OUT	STD_LOGIC;
	READY:			OUT	STD_LOGIC
);
END SHIFT_REGISTER;

ARCHITECTURE BEH OF SHIFT_REGISTER IS

	SIGNAL	DATA:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL	CONT: UNSIGNED(2 DOWNTO 0);
	
BEGIN	

DATAOUT	<=	DATA(0);
READY	<=	'1' WHEN (CONT="111") ELSE '0';

SR: PROCESS (cLK, RST, DATAIN, SHIFT_LOAD)
BEGIN
	IF(RST='1') THEN
		DATA<=(OTHERS=>'0');
		CONT<="000";
	ELSIF(RISING_EDGE(CLK)) THEN
		CASE SHIFT_LOAD IS
			WHEN "00" => NULL;
			WHEN "01" =>
				DATA	<=	STD_LOGIC_VECTOR(UNSIGNED(DATA) SRL 1);
				CONT<=CONT+1;
			WHEN OTHERS	=>
				DATA <= DATAIN;
				CONT<="000";
		END CASE;
	END IF;
END PROCESS;

END BEH;
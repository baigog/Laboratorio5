library ieee; 
use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;

--9600, 4800, 38400, 115200

--1- “Laboratorio 4: Completado por <Nombre_del_Alumno>”  
--2- “Curso 1er Escuela SE” 
--3- “<frase_a_eleccion_del_alumno>” 
--4- “<frase_a_eleccion_del_alumno>
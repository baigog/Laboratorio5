library ieee; 
use ieee.std_logic_1164.all;

ENTITY RS232_RX_FSM IS
	PORT(
		CLK:			IN	STD_LOGIC;
		RST:			IN	STD_LOGIC;
		TX:			IN	STD_LOGIC;
		PARITY_ERR:	IN	STD_LOGIC;
		
		SHIFT:			OUT	STD_LOGIC;
		DATA_OK:			OUT	STD_LOGIC;
		PARITY_CHECK:	OUT	STD_LOGIC
		);
END RS232_RX_FSM;

ARCHITECTURE BEH OF RS232_RX_FSM

SIGNAL CONT:	UNSIGNED(2 DOWNTO 0);
TYPE STATE IS (IDLE, START, DATA, PARITY, STOP);
SIGNAL CS, NS: STATE;
BEGIN

NEXT_STATE:	PROCESS (CS, TX, PARITY_ERR)
BEGIN
	CASE CS IS
		WHEN IDLE =>
			IF (TX=0) THEN
				NS <= START;
			ELSE
				NS <= IDLE;
			END IF;
		WHEN START => NS <= DATA;
		WHEN DATA =>
			IF (CONT = "111") THEN
				NS <= PARITY;
			ELSE
				NS <= DATA;
			END IF;
		WHEN PARITY => NS <= STOP;
		WHEN STOP =>
			IF(TX=1) THEN
				NS <= IDLE;
			ELSE
				NS <= STOP;
			END IF;
		WHEN OTHERS => NS <= IDLE;
	END CASE;
END PROCESS;

CURRENT_STATE: PROCESS (CLK, RST)
BEGIN
	IF(RST=1) THEN
		CS <= IDLE;
	ELSIF(RISING_EDGE(CLK)) THEN
		CS <= NS;
	END IF;
END PROCESS;

END BEH;
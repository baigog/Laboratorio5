library ieee; 
use ieee.std_logic_1164.all;

ENTITY LCD_CONTR_TB IS
END LCD_CONTR_TB;

ARCHITECTURE TB OF LCD_CONTR_TB IS

COMPONENT LCD_CONTR IS
	PORT(
			CLK:	IN STD_LOGIC	:= '0';		--RELOJ
			DATAIN:	IN	STD_LOGIC_VECTOR(7 DOWNTO 0)	:= (OTHERS=>'0');
			CLR:	IN STD_LOGIC	:= '0';
			WR:	IN STD_LOGIC	:= '0';
			RST:	IN STD_LOGIC	:= '0';
			
			EN:	OUT	STD_LOGIC;
			RWOUT:	OUT	STD_LOGIC;
			RS:	OUT	STD_LOGIC;
			LCD_ON:	OUT STD_LOGIC;
			BUSY:	OUT	STD_LOGIC;
			BL_ON:		OUT	STD_LOGIC;
			DATA:	INOUT	STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
END COMPONENT;

SIGNAL CLK, CLR,WR,RST:	STD_LOGIC:='0';	--ENTRADAS
SIGNAL DATAIN: STD_LOGIC_VECTOR(7 DOWNTO 0):= (OTHERS=>'0');
SIGNAL EN,RWOUT,RS,LCD_ON,BL_ON, BUSY:	STD_LOGIC;					--SALIDAS
SIGNAL DATA:	STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA_TX:	STD_LOGIC_VECTOR(7 DOWNTO 0)	:=	 (OTHERS=>'0');

BEGIN

LCD1: LCD_CONTR	PORT MAP(CLK=>CLK,DATAIN=>DATAIN,CLR=>CLR,WR=>wR, RST=>RST, 
									EN=>EN, RWOUT=>RWOUT, RS=>RS, LCD_ON=>LCD_ON, BL_ON=>BL_ON,
									BUSY=>BUSY, DATA=>DATA);

CLK	<=	NOT(CLK) AFTER 10ns;
DATA<=DATA_TX WHEN (RWOUT='1') ELSE (OTHERS=>'Z');

APLICA_ENTRADAS: PROCESS
BEGIN
	RST<='1';
	WAIT UNTIL RISING_EDGE(CLK);
	RST<='0';
	WAIT UNTIL FALLING_EDGE(BUSY);		--ESPERA HASTA FIN DE INICIALIZACION
	assert(false) report "INICIALIZACiON FINALIZADA" severity note;
	--FALTA PRUEBA DE ESCRITURA DE DATOS
	assert(false) report "FIN" severity failure;
END PROCESS;
END TB;
library ieee; 
use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;

--9600, 4800, 38400, 115200

ENTITY LABORATORIO5 IS
	PORT(
	
	);
END LABORATORIO5;


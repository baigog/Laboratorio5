library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY SHIFT_REGISTER_RX IS
PORT(
	CLK:				IN		STD_LOGIC;
	RST:				IN		STD_LOGIC;
	DATAIN:			IN		STD_LOGIC;
	SHIFT:			IN		STD_LOGIC;
	PARITY_OUT:		OUT	STD_LOGIC;
	DATAOUT:			OUT	STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END SHIFT_REGISTER_RX;

ARCHITECTURE BEH OF SHIFT_REGISTER_RX IS
SIGNAL	DATA:	STD_LOGIC_VECTOR(8 DOWNTO 0);
	
BEGIN
DATAOUT<=DATA(7 DOWNTO 0);
PARITY_OUT<=DATA(8);
SR: PROCESS (cLK, RST, SHIFT)
BEGIN
	IF(RST='1') THEN
		DATA<=(OTHERS=>'0');
	ELSIF(RISING_EDGE(CLK)) THEN
		IF (SHIFT='1') THEN
				DATA	<=	STD_LOGIC_VECTOR(UNSIGNED(DATA) SRL 1);
				DATA(8)	<= DATAIN;
		END IF;
	END IF;
END PROCESS;
END BEH;